module Top_proj (
    GPIO_LED1, //SINALIZAÇÃO START
    GPIO_LED2, //SINALIZAÇÃO START
    PMDO1_P7, //SCLK
    PMDO1_P8, //MOSI
    PMDO1_P9, //CS1
    PMDO1_P10, //CS2
    PMDO2_P1, //DHT
    PMDO2_P2, // DHT ERROR
    PMDO2_P3, // DEBUG
    CLK50MHZ //CLOCK PRINCIPAL
);

input CLK50MHZ;

output PMDO1_P7, PMDO1_P8, PMDO1_P9, PMDO1_P10, PMDO2_P2, GPIO_LED1, GPIO_LED2, PMDO2_P3; //SAÍDA PMOD
inout PMDO2_P1;

// wires para dht11
wire EN_DHT11,RST_DHT11, DHT_DATA, CRC_DHT, WAIT_DHT11, ERROR_DHT11;
wire [0:7] HUM_INT, HUM_FLOAT, TEMP_INT, TEMP_FLOAT;
reg EN_DHT11_REG, RST_DHT11_REG;
reg STARTED;
reg EN_DHT11_REG_START, RST_DHT11_REG_START;

assign PMDO2_P2 = ERROR_DHT11
//mULTIPLEXA A SAIDA ENTRE FSM START E PRICNIPAL
assign EN_DHT11 = STARTED ? EN_DHT11_REG: EN_DHT11_REG_START;
assign RST_DHT11 = STARTED ? RST_DHT11_REG: RST_DHT11_REG_START;

DHT11 DHT11(
    .CLK(BUFF50MHZ), // CLOCK PRICNIPAL
    .EN(EN_DHT11),
    .RST(RST_DHT11),
    .DHT_DATA(PMDO2_P1),
    .HUM_INT(HUM_INT),
    .HUM_FLOAT(HUM_FLOAT),
    .TEMP_INT(TEMP_INT),
    .TEMP_FLOAT(TEMP_FLOAT),
    .CRC(CRC_DHT),
    .WAIT(WAIT_DHT11),
    .error(ERROR_DHT11),
    .DEBUG(PMDO2_P3)

);
    
endmodule
